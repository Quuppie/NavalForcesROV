TRIODE PLATE CHARACTERISTIC CURVES
.DC LIN V_P 0 400 4    ; V_P IS THE SUPPLY VOLTAGE.  I(VP) IS OUTPUT.
V_P 101 0 200  ; PLATE VOLTAGE
VP 101 102 0   ; DUMMY VOLTAGE SOURCE FOR POSITIVE PLATE CURRENT PLOT.
VG 1 0 -1      ; GRID VOLTAGE.
R1 0 1 1G      ; ASSURES THAT GRID IS NOT FLOATING.

* X1 102 1 0 12AX7  ; P G C
* .STEP LIN VG 0 -4 .5    ; FOR 12AX7
X1 102 1 0 12AT7  ; P G C
.STEP LIN VG 0 -4 .5    ; FOR 12AT7
* X1 102 1 0 12AU7  ; P G C
* .STEP LIN VG 0 -20 4    ; FOR 12AU7
* X1 102 1 0 6DJ8   ; P G C
* .STEP LIN VG 0 -4 .5    ; FOR 6DJ8

.LIB C:\PSPICE\WORK\TUBE.LIB
.PROBE I(VG) I(VP)
.OPTIONS NOPAGE

* OLD TUBE MODELS FOLLOW FOR REFERENCE.

.SUBCKT TRIODE_12AX7 1 3 4  ; P G C
* 1 is plate; 3 is grid; 4 is cathode.  (2 is near plate.)
G1 2 4 VALUE={(EXP(1.5*(LOG((V(2,4)/93)+V(3,4)))))/680} ; S. REYNOLDS MOD.
C1 3 4 1.6P
C2 3 1 1.7P
C3 1 4 0.46P
R1 3 5 5000
D1 1 2 DX
D2 4 2 DX2
D3 5 4 DX
.MODEL DX D(IS=1P RS=1)
.MODEL DX2 D(IS=1N RS=1)
.ENDS

.SUBCKT TRIODE_12AU7 1 3 4  ; OLD MODEL
* 1 is plate; 3 is grid; 4 is cathode.  (2 is near plate.)
* G1 2 4 VALUE={(EXP(1.5*(LOG((V(2,4)/18)+V(3,4)))))/1151}
G1 2 4 VALUE=
+{EXP(PWR(V(2,4)/90*LOG(1+EXP(90*(1/20+V(3,4)/V(2,4))))),1.4)/790}
*    1   2 3   2       3     4   5      6   5  6   54321    0
C1 3 4 1.6P
C2 3 1 1.5P
C3 1 4 0.5P
R1 3 5 500
D1 1 2 DX
D2 4 2 DX2
D3 5 4 DX
.MODEL DX D(IS=1P RS=1)
.MODEL DX2 D(IS=1N RS=1)
.ENDS

.SUBCKT TETRODE_6L6 1 6 3 4  ; P G2 G1 C
G1 2 4 VALUE={((EXP(1.5*(LOG((V(6,4)/8)+V(3,4)))))/1455)*ATAN(V(2,4)/10)}
G2 6 4 VALUE={(EXP(1.5*(LOG((V(6,4)/8)+V(3,4)))))/9270}
C1 3 4 10P
C2 3 1 0.6P
C3 1 4 6.5P
R2 2 4 100K
D1 1 2 DX
D2 4 2 DX2
.MODEL DX D(IS=1P RS=1)
.MODEL DX2 D(IS=1N RS=1)
.ENDS

.SUBCKT TETRODE_6550 1 6 3 4  ; P G2 G1 C
G1 2 4 VALUE={((EXP(1.5*(LOG((V(6,4)/6.7)+V(3,4)))))/1455)*ATAN(V(2,4)/10)}
G2 6 4 VALUE={(EXP(1.5*(LOG((V(6,4)/6.7)+V(3,4)))))/9270}
C1 3 4 10P
C2 3 1 0.6P
C3 1 4 6.5P
R2 2 4 100K
D1 1 2 DX
D2 4 2 DX2
.MODEL DX D(IS=1P RS=1)
.MODEL DX2 D(IS=1N RS=1)
.ENDS

.END
